library verilog;
use verilog.vl_types.all;
entity comperator_vlg_vec_tst is
end comperator_vlg_vec_tst;
